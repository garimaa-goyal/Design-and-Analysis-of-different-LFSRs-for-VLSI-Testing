module lfsr_4bit_and_gate (   input clk,  input rst, output reg [3:0] q, output out, e,f);
reg [3:0] reg_q;
wire [3:0] q_wires;
wire e, f;

always @(posedge clk or posedge rst) begin
    if (rst) begin
        reg_q <= 4'b0001;
    end
     else begin
        if(reg_q[0] == 1'b0)
 begin
            reg_q = { reg_q[2], reg_q[3], reg_q[1], reg_q[0]}; // use blocking assignment
          reg_q <= {reg_q[0], reg_q[3] ^ reg_q[0],reg_q[2], reg_q[1]};
            q <= reg_q;
        end 
else 
begin
             reg_q <= {reg_q[0], reg_q[3] ^ reg_q[0],reg_q[2], reg_q[1]};
            q <= reg_q;
        end   
    end
end

assign q_wires = q;
assign e = ~(q_wires[3] & q_wires[2]);
assign f = ~(q_wires[1] | q_wires[0]);
and( out, e, f);

endmodule
